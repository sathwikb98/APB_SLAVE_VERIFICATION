`define ADDR_WIDTH 32      // Address bus width
`define DATA_WIDTH 32     // Data bus width
`define MEM_DEPTH 256     // Memory depth (number of locations)
